module baseline_test(
						clk_in         ,
						reset_in
					);



endmodule
